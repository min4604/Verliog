library verilog;
use verilog.vl_types.all;
entity and_not_or_vlg_check_tst is
    port(
        D               : in     vl_logic;
        E               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end and_not_or_vlg_check_tst;
