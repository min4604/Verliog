library verilog;
use verilog.vl_types.all;
entity and_not_or_vlg_vec_tst is
end and_not_or_vlg_vec_tst;
